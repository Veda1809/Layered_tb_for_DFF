interface intf(input bit clk);
  
  logic D;
  logic reset;
  logic Q;
  
endinterface
